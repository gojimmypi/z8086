(* blackbox *)
module OBUFDS (
    input  wire I,
    output wire O,
    output wire OB
);
endmodule

(* blackbox *)
module ODDRX1F (
    input  wire D0,
    input  wire D1,
    input  wire SCLK,
    input  wire RST,
    output wire Q
);
endmodule
