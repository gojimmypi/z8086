(* blackbox *)
module pll27 (
    input  wire clkin,
    output wire clkout0,
    input  wire mdclk
);
endmodule

(* blackbox *)
module pll74 (
    input  wire clkin,
    output wire clkout0,
    output wire clkout1,
    input  wire mdclk
);
endmodule
